module top_module ( input a, input b, output out );
    mod_a test1 (.out(out), .in2(b), .in1(a));
    
endmodule
