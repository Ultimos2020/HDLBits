module top_module( input in, output out );
wire t;
    assign t = in;
    assign out = t;
    
endmodule
